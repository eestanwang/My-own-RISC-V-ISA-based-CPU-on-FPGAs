module and_3 (
    input  a,
    output b
);
  and_2 and_2_inst (
      .a(a),
      .b(a),
      .c(b)
  );

endmodule  //and_3
