module and_2 (
    input  a,
    input  b,
    output c
);

  assign c = a & b;
endmodule  //and_2
